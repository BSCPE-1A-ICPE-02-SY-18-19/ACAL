CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 110 10
176 80 1278 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 218 152 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3751 0 0
2
43530.4 0
0
6 74LS48
188 851 177 0 14 29
0 3 6 5 4 17 18 8 9 10
11 12 13 14 19
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4292 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 963 73 0 18 19
10 14 13 12 11 10 9 8 20 21
1 0 0 1 0 1 1 2 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6118 0 0
2
43530.4 1
0
9 2-In AND~
219 622 112 0 3 22
0 7 6 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
34 0 0
2
43530.4 2
0
9 2-In AND~
219 484 111 0 3 22
0 4 5 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6357 0 0
2
43530.4 3
0
7 Pulser~
4 105 321 0 10 12
0 22 23 24 15 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
319 0 0
2
5.89883e-315 0
0
6 74112~
219 697 277 0 7 32
0 2 16 15 16 2 25 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3976 0 0
2
5.89883e-315 5.26354e-315
0
6 74112~
219 549 277 0 7 32
0 2 7 15 7 2 26 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7634 0 0
2
5.89883e-315 5.30499e-315
0
6 74112~
219 392 277 0 7 32
0 2 4 15 4 2 27 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
523 0 0
2
5.89883e-315 5.32571e-315
0
6 74112~
219 258 277 0 7 32
0 2 28 15 29 2 30 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6748 0 0
2
5.89883e-315 5.34643e-315
0
35
1 0 2 0 0 8192 0 1 0 0 23 4
218 164
218 184
258 184
258 189
7 1 3 0 0 8320 0 7 2 0 0 4
721 241
753 241
753 141
819 141
0 4 4 0 0 8320 0 0 2 25 0 3
330 241
330 168
819 168
0 3 5 0 0 12416 0 0 2 32 0 4
439 240
458 240
458 159
819 159
0 2 6 0 0 12416 0 0 2 31 0 4
590 241
621 241
621 150
819 150
0 0 2 0 0 4096 0 0 0 9 23 2
633 289
633 189
0 0 2 0 0 0 0 0 0 10 23 2
469 289
469 189
0 0 2 0 0 0 0 0 0 23 11 2
312 189
312 289
5 5 2 0 0 4096 0 8 7 0 0 2
549 289
697 289
5 5 2 0 0 4096 0 9 8 0 0 2
392 289
549 289
5 5 2 0 0 0 0 10 9 0 0 2
258 289
392 289
2 0 7 0 0 4096 0 8 0 0 13 2
525 241
505 241
4 3 7 0 0 8320 0 8 5 0 0 3
525 259
505 259
505 111
7 7 8 0 0 4224 0 2 3 0 0 3
883 141
978 141
978 109
8 6 9 0 0 4224 0 2 3 0 0 3
883 150
972 150
972 109
9 5 10 0 0 4224 0 2 3 0 0 3
883 159
966 159
966 109
10 4 11 0 0 4224 0 2 3 0 0 3
883 168
960 168
960 109
11 3 12 0 0 4224 0 2 3 0 0 3
883 177
954 177
954 109
12 2 13 0 0 8320 0 2 3 0 0 3
883 186
948 186
948 109
13 1 14 0 0 8320 0 2 3 0 0 3
883 195
942 195
942 109
1 0 2 0 0 0 0 8 0 0 23 2
549 214
549 189
1 0 2 0 0 0 0 9 0 0 23 2
392 214
392 189
1 1 2 0 0 8320 0 7 10 0 0 4
697 214
697 189
258 189
258 214
2 0 4 0 0 0 0 9 0 0 25 2
368 241
355 241
7 0 4 0 0 0 0 10 0 0 26 2
282 241
355 241
1 4 4 0 0 0 0 5 9 0 0 4
460 102
355 102
355 259
368 259
3 0 15 0 0 8192 0 10 0 0 35 3
228 250
206 250
206 321
3 1 7 0 0 0 0 5 4 0 0 3
505 111
505 103
598 103
2 0 16 0 0 4096 0 7 0 0 30 2
673 241
653 241
3 4 16 0 0 8320 0 4 7 0 0 4
643 112
653 112
653 259
673 259
7 2 6 0 0 0 0 8 4 0 0 4
573 241
590 241
590 121
598 121
2 7 5 0 0 0 0 5 9 0 0 4
460 120
439 120
439 241
416 241
3 0 15 0 0 0 0 8 0 0 35 3
519 250
487 250
487 321
3 0 15 0 0 0 0 9 0 0 35 3
362 250
340 250
340 321
4 3 15 0 0 4224 0 6 7 0 0 4
135 321
641 321
641 250
667 250
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
